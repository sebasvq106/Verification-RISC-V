`include "top_hvl.sv"
`include "interface.sv"
`include "riscv_item.sv"
`include "sequence.sv"
`include "driver.sv"
`include "monitor.sv"
`include "scoreboard.sv"
`include "coverage.sv"
`include "assertions.sv"
`include "agent.sv"
`include "env.sv"
`include "test_1.sv"
`include "test_r_type.sv"
`include "test_i_type.sv"
`include "test_load_type.sv"
`include "test_store_type.sv"
`include "test_lui_type.sv"
`include "test_reset.sv"
