interface intf_cnt(input tb_clk);
  
  logic reset;
  logic [31:0] tb_WB_Data;

endinterface
  
  