`include "../testbench/top_hvl.sv"
`include "../testbench/interface.sv"
`include "../testbench/riscv_item.sv"
`include "../testbench/sequence.sv"
`include "../testbench/driver.sv"
`include "../testbench/monitor.sv"
`include "../testbench/scoreboard.sv"
`include "../testbench/agent.sv"
`include "../testbench/env.sv"
`include "../testbench/test_1.sv"

