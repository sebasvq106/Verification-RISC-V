`include "top_hvl.sv"
`include "interface.sv"
`include "driver.sv"
`include "env.sv"
`include "test_1.sv"
