`include "../testbench/top_hvl.sv"
`include "../testbench/interface.sv"
`include "../testbench/riscv_item.sv"
`include "../testbench/sequence.sv"
`include "../testbench/driver.sv"
`include "../testbench/monitor.sv"
`include "../testbench/scoreboard.sv"
`include "../testbench/assertions.sv"
`include "../testbench/agent.sv"
`include "../testbench/env.sv"
`include "../testbench/test_1.sv"
`include "../testbench/test_load_type.sv"
`include "../testbench/test_store_type.sv"
`include "../testbench/test_lui_type.sv"
`include "../testbench/test_i_type.sv"
`include "../testbench/test_r_type.sv"
`include "../testbench/test_reset.sv"