class scoreboard;
  
 	logic [31:0] instruction_queue [$];

endclass