`include "../testbench/interface.sv"
`include "RISC_V.sv"
`include "top_hdl.sv"
