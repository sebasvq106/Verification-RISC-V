`include "RISC_V.sv"
`include "top_hdl.sv"