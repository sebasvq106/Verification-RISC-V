`include "RISC_V.sv"
